module Exnorgate (
input a,b,
output y
);
xnor (y,a,b);
endmodule
