module norgate (
input a,b,
output y
);
nor (y,a,b);
endmodule
