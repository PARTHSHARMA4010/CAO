module notgate (
input a,
output y
);
not (y,a);
endmodule
