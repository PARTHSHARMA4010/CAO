module andgate (
input a,b,
output y
);
and (y,a,b);
endmodule
