module orgate (
input a,b,
output y
);
or (y,a,b);
endmodule
