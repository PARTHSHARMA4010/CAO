module Exorgate (
input a,b,
output y
);
xor (y,a,b);
endmodule
