module Exnorgate_test;
reg a,b;
wire y;
Exnorgate uut(a,b,y);
initial begin 
$dumpfile("Exnorgate.vcd");
$dumpvars(0,Exnorgate_test);
a=0;b=0;
#10
a=0;b=1;
#10
a=1;b=0;
#10
a=1;b=1;
#10
$finish();
end
endmodule
